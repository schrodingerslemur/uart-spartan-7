��m o d u l e   t o p   (  
         / /   U A R T   i n t e r f a c e  
         i n p u t     l o g i c   b l e _ u a r t _ r x ,  
         i n p u t     l o g i c   C L O C K _ 1 0 0 ,  
         o u t p u t   l o g i c   b l e _ u a r t _ t x ,  
  
         / /   L E D s  
         o u t p u t   l o g i c   [ 1 5 : 0 ]   L E D ,  
  
         / /   B u t t o n s  
         i n p u t     l o g i c   [ 3 : 0 ]   B T N ,  
  
         / /   S w i t c h e s  
         i n p u t     l o g i c   [ 1 5 : 0 ]   S W ,  
  
         / /   A n o d e s   a n d   s e g m e n t s  
         o u t p u t   l o g i c   [ 3 : 0 ]   D 1 _ A N ,   D 2 _ A N ,  
         o u t p u t   l o g i c   [ 7 : 0 ]   D 1 _ S E G ,   D 2 _ S E G  
  
 ) ;  
  
     l o g i c   e n ;  
  
     / /   I n s t a n t i a t e   U A R T   m o d u l e  
     u a r t   # (  
         . B A U D _ R A T E       ( 1 1 5 _ 2 0 0 ) ,  
         . C L O C K _ F R E Q     ( 1 0 0 _ 0 0 0 _ 0 0 0 ) ,  
         . D A T A _ B I T S       ( 8 )  
     )   u a r t _ i n s t   (  
         . c l o c k             ( C L O C K _ 1 0 0 ) ,  
         . r e s e t             ( B T N [ 0 ] ) ,  
         . t x _ d a t a         ( S W [ 7 : 0 ] ) ,                     / /   E x a m p l e   d a t a   t o   s e n d  
         . t x _ s e n d         ( B T N [ 1 ] ) ,                   / /   S e n d   d a t a   o n   b u t t o n   p r e s s  
         . t x _ b u s y         ( ) ,                                 / /   U n u s e d   i n   t h i s   e x a m p l e  
         . r x _ d a t a         ( ) ,  
         . r x _ v a l i d       ( e n ) ,  
         . r x                   ( b l e _ u a r t _ r x ) ,  
         . t x                   ( b l u e _ u a r t _ t x )  
     ) ;  
  
         / /   R e g i s t e r  
         a l w a y s _ f f   @ ( p o s e d g e   C L O C K _ 1 0 0   o r   p o s e d g e   B T N [ 0 ] )   b e g i n  
                 i f   ( B T N [ 0 ] )   b e g i n  
                 L E D   < =   1 6 ' b 0 ;  
                 e n d   e l s e   i f   ( e n )   b e g i n  
                 L E D   < =   { 8 ' b 0 ,   u a r t _ i n s t . r x _ d a t a } ;   / /   D i s p l a y   r e c e i v e d   d a t a   o n   l o w e r   8   L E D s  
                 e n d  
         e n d  
  
 e n d m o d u l e :   t o p  
 